library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;

entity PhaseCalibration is
	generic (
		BOARD_ID : integer := 0
	);
	port (
		clk			  : in  std_logic;
		phase_in	 	  : in  std_logic_vector (6 downto 0);
		amplitude_in  : in  std_logic_vector (6 downto 0);
		color_in		  : in  std_logic_vector (26 downto 0);
		address_in	  : in  std_logic_vector (7 downto 0);
		phase_out	  : out std_logic_vector (6 downto 0);
		amplitude_out : out std_logic_vector (6 downto 0);
		color_out 	  : out std_logic_vector (26 downto 0)
	);
end PhaseCalibration;

architecture Behavioral of PhaseCalibration is

	subtype CALIB_PHASE is std_logic_vector(6 downto 0);
	type CALIBLATION_ROM is array (0 to 255) of CALIB_PHASE;
	constant calib_rom_0 : CALIBLATION_ROM := (
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000",
		"0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000", "0000000"
	);	
	constant calib_rom_1 : CALIBLATION_ROM := (
		"0110110","0111000","1111010","0101101","0110100","0110001","1110100","1101100","1110111","0110000","1110011","0110010","0101101","1110100","0110001","0101010",
		"0110111","0110001","0101111","0110100","0110010","0101110","0110011","0110110","0110110","0100111","0110100","1110110","0110010","0110100","0110001","1110001",
		"1110101","1111000","0110110","1110111","1110101","0110100","1110101","1110111","0110101","0110001","0110011","0110100","1110100","1110110","1111000","1110011",
		"0110011","0110011","0111000","0110100","0110100","0110011","1110110","1110011","0110010","0110011","0110100","0110101","1110110","1110010","0110101","1110100",
		"0111011","1110010","0110100","0110011","1110101","0001100","0110110","0110101","0110101","0110011","0110010","0110101","0110011","0110100","1110011","0111000",
		"1110101","1110111","0110010","0110010","0110101","1110111","0110110","0110101","1110101","0110111","0110100","0110011","1111000","0110111","1110101","1110010",
		"0111000","0110100","0110100","0110000","1110100","1110000","0110011","0110111","0111000","1110100","0110110","1110110","1110111","1110011","1110111","1110011",
		"0110111","1110011","1110100","0110110","0111000","0111010","0110110","0110110","1110100","0101111","0110010","1110100","1110111","0110100","1110110","1110011",
		"0110101","0111000","1110010","0110001","0111011","0110011","1110010","1110110","1110100","0110010","1111000","0110110","0110100","1110101","0110011","0110101",
		"0110011","0110110","0110010","1111001","0110100","0110001","0110001","1110001","0110101","1110100","0110101","0110100","0110100","1110111","1110101","0110000",
		"0110000","0110110","0110010","0110011","0101111","1110110","0110111","1101100","0110110","1110110","1110011","1110100","1111001","0110110","1110100","0101111",
		"1110110","0110101","1110101","0110111","0110101","0111010","0110101","0110101","0111000","0110111","0110011","0111000","1110001","1110101","1110111","1110011",
		"0110110","0101110","0110010","1110101","1110001","0110100","0110101","0111001","0110100","1111000","1111100","1110110","0111001","0110100","0101111","1110101",
		"1110101","0110110","1110110","0110100","1111011","0110111","0110100","1111000","1110101","0110110","1110011","0110010","1110000","1110101","1101110","0110001",
		"0110100","1110111","0110100","0110001","0110100","0110110","1111001","1110110","0110101","0110000","1110100","1111000","1110011","0110100","0110111","1110010",
		"0110011","1110101","1111100","0110101","1110110","1101111","0111010","0110100","1110111","1110000","0101011","0110011","0110110","1110100","1110100","1110110"
	);
	constant calib_rom_2 : CALIBLATION_ROM := (
		"0010000","1010000","0001010","0010000","1010101","0001110","0010101","1001100","0000000","1001110","0001110","0010101","1010000","0001010","1010001","0001110",
		"1001100","1010000","0001100","1010001","0010011","0001110","1001010","0000111","1010001","0010001","1001110","1001000","0001110","1000101","0000101","1001000",
		"1001110","1010001","1001110","0001100","0001110","1001110","1001010","1001010","1001110","1000111","1010000","0001010","0001000","1010001","1001100","0000111",
		"0010000","0000101","0001110","1001000","1010011","0001010","0001010","1001010","0001100","0001010","0000011","0001100","1001110","1001110","1010001","1001110",
		"0010101","0010101","1001010","0001100","0010001","1010000","1001010","0010000","1010000","0010000","1000001","1001010","1010000","0000111","0001010","1010000",
		"0010000","0000111","0001010","0000111","1001110","1010000","1000101","0010000","1010000","0010001","0000101","1001010","0000011","1010001","0001110","1010000",
		"1010001","0010001","1010000","1001110","1001000","1001000","0001110","1010001","0010000","0001010","1010001","1001110","1001100","1010000","0000101","0001110",
		"1010101","0001110","0010001","0001010","0001110","0001000","1001110","1010001","1001100","0001010","1010001","0010000","0010011","0010001","0010101","0001110",
		"0011010","0001010","1000101","1001010","1001010","0001100","1011000","0001110","0010011","1001010","0010001","0110001","0001010","1010000","0001100","0001110",
		"0010001","1001010","1001010","1011010","1001000","0001010","0001010","0001010","1001110","1010001","1001110","1011100","0010000","1010101","0010001","0010001",
		"0000101","1000101","1001110","1010000","0001010","1010101","1010101","1001110","0011000","0001010","1001010","1001110","1010101","0000111","0010011","0001010",
		"0001100","0010000","1010001","0001110","1010000","0010001","1001100","0001000","0000001","0010001","1010001","1001110","0001010","1001110","0010001","1010001",
		"1010101","1011100","1010000","1001010","0001100","1001110","0001100","0010001","0001010","1001100","0001110","0001010","1001110","0011110","0010001","1010001",
		"0001100","1011010","0001110","1010001","1000101","1000111","1010000","1010001","0001110","1010000","1001010","0011010","1001000","1010000","1001010","1010001",
		"0001110","0001010","1010001","0000101","1000011","0001110","1001110","0001000","0010000","1001010","0001110","0010001","1010001","0010011","1001010","1010101",
		"1010000","0011000","0010001","1010001","0001100","1001110","0001000","0011000","1001010","1001010","1010001","1010001","0010000","1001010","1001010","1001110"
	);
	constant calib_rom_3 : CALIBLATION_ROM := (
		"1110100","0110101","0111000","0110111","0110010","0110010","0110001","1110100","0110011","0111001","1110110","1111000","1110110","0110010","1101111","0110001",
		"0110101","0110101","1110110","0110011","0111000","0110111","1110100","1111001","0110101","1110111","1110100","1111000","1110111","1110110","0110010","0111000",
		"1110011","0111000","0110100","0110101","1111001","0110111","0110011","0110110","0110101","1110100","0110110","1110110","0110110","0110100","0110010","1110100",
		"1110011","1110100","0001100","0110100","0110011","1110111","0110100","1110111","1110100","0110010","1111000","1111000","1110011","1111000","0110101","0110001",
		"0110101","1110110","1110001","1110100","0110101","1110111","1110100","0111010","1110100","0110101","0111000","0110101","1110110","0110100","0111000","0110101",
		"0110101","1110111","0110101","1110010","0110001","1111111","1110010","1110111","0110100","1110101","0110110","0111000","1110000","0110010","1110100","0110010",
		"1110110","1111000","0110001","0110101","1110111","0110000","1110110","1111001","0110011","1110010","0110101","0110010","1110101","1110111","1110100","0110111",
		"0111011","0110010","1110110","0111001","0110101","0110110","0111001","0111000","1110110","0110101","1110101","1111100","1111000","0110001","1110100","0110101",
		"1110111","0110101","0110010","0111000","0111001","0111010","1110101","0111000","1110111","1111100","0111001","0110111","1110100","1110110","1110110","0111000",
		"0110011","0111000","0110101","0110100","0111001","1110100","0110100","0110110","0110100","1110111","0000111","1110100","1110011","0110010","0110001","1110111",
		"0110001","1111000","0110011","1110001","0110111","0110100","0111000","0101101","0110100","0110110","0111100","1111100","0111001","0110101","0110101","0110011",
		"0111100","0110101","0110010","1110101","0110011","1110011","1111001","0110111","0110101","0110001","1110101","1110011","0110111","0110110","1111000","1110101",
		"1110100","0110011","0110011","0110110","0110100","0110100","1110111","1110110","1110010","0110110","1110101","0110101","0110101","1110100","1110101","0110100",
		"1111010","0110110","1110011","1110111","0101111","1110111","1110001","0110111","1110100","1111001","1110110","0110111","1110110","1110100","0110010","0111011",
		"0110110","0110100","1110011","0110110","0110110","0110111","0111001","1110010","0110111","1110111","1110111","0110010","0110111","0110011","1110011","1111000",
		"0110101","0110100","0110001","0110110","1110100","1111100","0111000","1110100","0110110","0110011","1110010","1110000","1110111","0110001","0110111","1110100"
	);
	constant calib_rom_4 : CALIBLATION_ROM := (
		"1110111","0111010","1110001","0110110","0110010","0110100","0110101","1111001","0110011","1110010","0110101","0111010","0110101","1110011","1110101","1111010",
		"0110101","0111100","1111001","0110101","1111000","0111100","1110111","1110110","1101110","1111010","0000000","1110111","1110011","0110000","1111010","1110110",
		"0110110","0111001","1110100","1111010","1111000","1111000","0111010","1111000","0110111","0111000","0110000","0110011","0110101","0110011","1111000","1110111",
		"0110011","1110110","1110111","0111011","1110101","0111001","1111000","1111001","1111000","0110110","0110110","0110011","0110111","1110111","0111001","0110001",
		"1110110","0110111","1110011","1110111","1110101","1110101","0111001","0110101","0110110","0110011","1110100","1110100","0110110","1111011","0111000","0110010",
		"1110101","1110101","1110110","0110111","0110001","1111000","0110110","1110111","1110110","1110100","1110101","0110110","1110101","1110010","0110101","1110101",
		"0110110","0110101","1110110","0110001","0110100","1110100","1110111","1110111","1110111","1111000","1110010","1110011","0110101","0111010","1110101","0110000",
		"1110110","1111000","1111000","1110110","1110111","0110111","0110101","1110101","0110110","0110101","1110011","0110011","0110111","0110100","1110010","1110001",
		"0110111","1110101","0111011","0111000","1110110","1110110","1110111","1110111","1110110","0110001","0111001","1110111","1111011","0110110","1110111","1110110",
		"0111000","0110011","1110111","1110111","1111001","0111001","1110100","1110100","1110110","0110110","0110011","1110111","1110011","0110101","1110110","1110111",
		"1110111","0110111","1111000","0110100","1111000","1111000","1110101","1110011","1110111","0110011","1110101","1110001","0110101","0110101","0110111","0110001",
		"1111000","0110001","1110101","1110100","0110100","0110011","1110111","1110101","0110101","0111000","1110010","1111000","0110100","1111000","0110110","0110110",
		"1110100","0110111","1110110","0110010","1110110","1110111","1110001","0110101","0110001","1110100","0110101","1110111","0110111","0111000","0111000","0110111",
		"0110100","0111000","0111100","1110100","1110011","0110110","1110100","1110110","0111000","1110100","1110110","1110110","0110110","1111000","0110111","0110100",
		"1110100","1110110","1110101","0110110","1110111","1110110","1110111","0110100","1110001","0110101","0110011","1110110","1110010","1110100","0110100","1110010",
		"0110011","1110001","1110110","0110100","1110111","0110110","1110110","0110101","1110100","1111001","1110111","1110111","1110100","1110000","1110011","1110011"
	);
	constant calib_rom_5 : CALIBLATION_ROM := (
		"1110011","1110011","1110110","1110101","0111100","1110100","0110110","1110011","0110100","0111000","1101010","1110011","0110111","1111000","1110101","0110000",
		"0111011","1110111","0110111","1110110","1110100","1110111","0111000","1111011","0111000","1110011","0111001","1110110","0111001","0110101","0111001","0110011",
		"0111000","0110101","1110111","1110111","1110100","1110010","0111001","0110100","0110011","1110111","0110010","0110100","1110111","0110110","0110101","0110100",
		"0110110","1000000","0111000","0110101","0110111","0110101","0111000","1110100","0110100","0110110","0111000","0111000","0111000","1110101","0110101","1110111",
		"1110111","0110010","0110110","0111000","1110100","1110111","1110111","1110011","1111000","1110101","1101100","1110011","1110010","0110110","1111010","1110111",
		"0110101","0110110","1111010","1110110","0110100","1110101","1110100","1111010","1111011","0110110","1111000","0110111","1110110","0110110","1110010","0110101",
		"0110101","0110011","1110110","0110110","1110100","0110111","1110110","0110001","1110110","0110101","0110101","0110111","1110110","1110110","1110011","1110011",
		"1110100","0111000","0110110","0110111","0110101","0110110","1111001","0110110","0110011","0110100","0110110","0110011","1110101","1110010","1110110","0110101",
		"1111100","0110111","1110111","0111000","1110101","0110111","0110011","0110100","0110101","1110111","1110001","1110110","0110100","0110100","1111011","1111000",
		"1111001","1110100","1110001","1110011","0110110","1110011","0110100","0110111","1110011","1110110","1110100","1111000","1110101","0111000","0110010","1110101",
		"1110110","1110101","1110011","1110111","1110100","1110101","1111001","1110111","0110101","0110101","0110110","0110110","0110010","0110100","0110010","1110101",
		"0110111","1110010","0111001","1110111","1110110","0110001","0110100","1110100","0111001","1110100","1110100","0110110","1110100","1110111","1111001","0110100",
		"1110100","0110101","0110101","0111001","1110100","0110100","1111001","0110100","0110101","0110010","1110011","1110011","1110101","0110011","0110100","1111011",
		"1110101","0110100","0110100","0110111","0110100","1110101","0111000","1110101","1110110","0111011","1110101","1110111","1110110","1110101","1110011","0110001",
		"0110010","0110100","0110100","1110101","0110100","0111000","0110101","1110110","0110101","1110001","0110101","0101110","1110011","1110100","1110011","1110100",
		"1110111","1110100","0110011","0111000","0100110","0110011","0110000","0110101","0111001","1110100","0110011","0110001","1110100","1101001","1110101","0110101"
	);
	constant calib_rom_6 : CALIBLATION_ROM := (
		"0110000","0111010","0110011","0110101","0110010","1110001","0110011","0110010","0110000","0110010","1110010","1110111","1110100","1110010","0101111","0110001",
		"0110011","1110011","0110011","1110101","1110100","0110010","0110010","0110011","0110001","0110000","1110010","1110010","1110011","1110100","1110011","1110011",
		"1110011","0110010","1110000","1110010","1110110","0110010","1110010","0110100","1110111","0110001","0110100","0110011","0110100","0111001","1110100","1110001",
		"1110100","0110010","0110001","0110010","1110101","0110101","1110011","0110010","1110011","0110010","0110010","1110011","1110010","1110011","0110011","1110110",
		"1110011","1110000","0110100","0110110","0110110","0110001","0110110","0110110","0110000","1111001","1110011","1110010","1110011","0110010","1110010","1110101",
		"0110010","1110000","0110101","0110110","0110110","0110001","0110101","0110011","0110000","1110111","1110010","1110000","1110011","0110001","1110011","1110101",
		"0110011","1110010","0110101","0110010","0110100","0110000","0110000","1110110","1110100","0110100","1110100","0110010","0110010","1110100","0110110","1110111",
		"0110010","0110010","0110011","0110001","1110001","0110010","0110100","0110011","1110100","0110010","0110011","1110000","1110000","1110010","1110001","0110110",
		"0110000","1110100","1110001","1110101","1110110","0110001","1110100","1110011","1110110","1110100","1110011","1110010","0110100","1110101","0110011","1110101",
		"1110101","0110101","1110011","1110011","0110011","1110101","0110100","1110010","0110010","0110100","1110010","1110011","1110001","1110001","1110011","0110001",
		"1110100","0110100","1110100","1110000","1110001","1110101","0110100","1110011","0110011","1110010","0110101","1110010","1110011","0110010","0110011","1110101",
		"1110011","0110110","1110011","0110101","0110010","1110100","1110101","0110011","1110100","1110001","0110001","0110100","1110011","1101111","0110000","0110010",
		"1110000","1110100","0110101","1110010","1110011","0110100","1110010","0110100","1110001","0110010","0110001","0110010","1110110","1110000","0110011","0110100",
		"0110100","1110001","1110111","0110000","0110100","0110000","1110011","0110011","1110100","0110000","1110001","0110010","1110101","0110011","1110011","0110100",
		"1110111","1110010","0101110","0101110","0110100","0110010","1110011","0110011","0110001","0110011","1110011","0110100","0110001","0110110","0110011","1110100",
		"0110010","1110000","0110011","1110001","1110110","0110001","0110001","1110100","1110101","1110101","0110010","1110000","1101110","0110010","0110001","1110010"
	);
	constant calib_rom_7 : CALIBLATION_ROM := (
		"1001010","0001000","0000111","1000011","1000011","0000011","1001010","0000000","0000000","1000001","1000011","1000001","0000000","0000000","1000111","1001000",
		"1000011","0001000","0000011","1000011","1111110","0010001","0001000","0000011","0000000","1000101","1000111","1000000","0000000","0000001","1000111","1000111",
		"1000001","0001010","1000000","1111110","1000001","0000000","0000111","1000011","1000001","0111110","1000001","1000000","0000011","0000001","0000101","1001000",
		"1000111","1000011","0000101","1000001","0000000","1000011","0111100","0000101","0111100","0000111","1000011","0000011","0000011","1111110","1000001","1001110",
		"0000000","0001000","1000001","0111110","0000011","0000111","0000101","0000111","0000001","0001000","1000011","0000001","1000111","1000000","1000111","0001100",
		"1111100","0000101","0111100","1000000","1000001","1000001","0001010","0000000","1001000","1000011","0000101","0000000","1000011","1001010","0000111","1001010",
		"0111100","0000011","1000111","1000011","1000000","0000000","0000011","0000001","0000000","1000111","1000111","1000111","0111100","0000011","1011000","0001010",
		"0000000","0000101","0001110","1000011","1000000","0000101","0111110","1000001","1001010","0000111","0000101","1000111","1000011","0001110","0000011","0001010",
		"1000001","1000011","1000111","1000011","0000111","0000101","0000111","0000011","0000001","1000111","1001010","1000011","0000001","0000111","1000111","1001000",
		"1000111","0000011","0000000","1111100","0000000","1000011","0000011","1000111","1000011","1000011","1001100","0001000","1111100","0000000","1000001","0001000",
		"0000000","0000011","1111100","1000011","0000011","1001110","0001100","0000011","0001000","0000011","0000111","1000001","1000111","1000111","1000111","1000101",
		"1000000","0000011","0000111","1000101","0111110","1000111","0001010","1000000","0000101","1000011","0000111","1000101","0000111","0001010","1001010","1000111",
		"1000000","0000011","1010000","0000011","1000101","0000000","0000111","0000111","0000000","0000001","0000101","0000101","1000000","1001010","0001010","1001100",
		"1000001","1000111","1000111","0000000","0000001","0111110","0000101","0000001","0000011","0001010","0000111","1000011","1010000","0001010","1000111","0000111",
		"0000111","1010011","0000011","1000001","0000001","0000000","0000000","1000000","0000011","0000011","0000111","0000000","1000111","1001100","0001010","0000001",
		"0001010","0001110","0000011","0000011","1001000","1000001","0000001","0000011","1000011","1001010","0000111","1001100","0000111","0001010","1001110","0001100"
	);
	constant calib_rom_8 : CALIBLATION_ROM := (
		"1110011","1110111","1110101","1110011","1110101","1110101","0110011","1110101","0111000","0110111","0110101","1000001","1100111","0000011","0001100","0000111",
		"0110101","0110101","0110101","0110111","1111000","1110001","0110001","0110101","1111000","1111000","0111000","0111100","1011100","0100001","1011100","1011100",
		"0110000","0110101","1110111","1110101","1110011","0110001","1110011","0111000","1110101","0111000","0110111","0111010","1000001","1111000","1100111","1010101",
		"1110001","1111000","0110011","1110000","0110011","1110011","0110101","0110111","0111000","0110101","1111000","0010101","1000111","1110000","0100000","1111110",
		"1111100","0110111","1110001","1101110","0110101","1110011","1110001","1011000","0111000","1111000","0111000","1000001","1101010","1010011","0111000","0011010",
		"0110000","1110111","0010001","0110001","0110101","1110011","0110101","0111000","1111000","0011000","0111000","1111100","0101110","0010101","1110001","1011000",
		"1110001","1110101","0110001","0110001","0111000","0110101","1110101","1110111","1111000","0110111","1110111","0000111","0111110","0110000","0011100","1000001",
		"0110011","0111000","1110001","1110001","1110101","0110001","1110101","1111000","1111100","0000000","1111010","1101010","1101110","0110001","0101010","1010101",
		"1110101","0110101","1110101","0110001","1110000","0111000","1110101","0111000","1111000","0110111","1111000","1111000","1001110","1011010","1011000","1010101",
		"1110101","1110101","1110001","0110101","0110011","0110011","1110101","1111000","0111000","1110111","0000000","0111010","0100101","0111100","0000101","0000111",
		"0101110","0110001","1110101","1110101","1110101","0110011","1110001","1111010","0111000","0110111","0111100","1110001","1100000","0001000","0100000","0101000",
		"0111000","0110101","1110001","1110011","1110101","1110011","1110101","0111000","1111100","0001010","0111100","0100011","0100101","1001110","1101010","1111000",
		"0110011","0010000","0110001","0110101","1001010","0110001","1111000","1110111","1111100","0111010","0111000","1010001","0011000","0001000","0110001","0010000",
		"0110011","0110000","0110001","1110011","0110001","1110101","1110101","0110011","1111000","1000001","1111000","0111110","0001010","0000011","1110001","1010011",
		"0110000","0110001","0110011","1110011","1110101","1110001","1110001","1110111","0110111","0110111","1111000","0101010","1111100","0111110","0110001","1011000",
		"0110011","1110011","1110001","1110101","0110111","1111000","1110111","1110101","1111000","0111000","0111100","1010101","0101010","1110001","0101110","1011000"
	);
	
	
	signal original		  : std_logic_vector (7 downto 0) := (others => '0');
	signal calib_out  	  : std_logic_vector (6 downto 0) := (others => '0');
	signal amplitude_out_d : std_logic_vector (6 downto 0) := (others => '0');
	signal color_out_d	  : std_logic_vector (26 downto 0) := (others => '0');
	signal phase_out_s 	  : std_logic_vector (7 downto 0) := (others => '0');
	signal amplitude_out_s : std_logic_vector (6 downto 0) := (others => '0');
	signal color_out_s	  : std_logic_vector (26 downto 0) := (others => '0');

begin

	phase_out <= phase_out_s(6 downto 0);
	amplitude_out <= amplitude_out_s;
	color_out <= color_out_s;

	process (clk) begin
		if rising_edge(clk) then
			case BOARD_ID is
				when 0 => 
					calib_out <= calib_rom_0(CONV_INTEGER('0' & address_in));
				when 3 =>
					calib_out <= calib_rom_3(CONV_INTEGER('0' & address_in));
				when 7 =>
					calib_out <= calib_rom_7(CONV_INTEGER('0' & address_in));				
				when others =>
					calib_out <= calib_rom_0(CONV_INTEGER('0' & address_in));
			end case;
					
			original <= ("0" & phase_in);
			phase_out_s <= original - ("0" & calib_out);
			
			amplitude_out_d <= amplitude_in;
			amplitude_out_s <= amplitude_out_d;
			color_out_d <= color_in;
			color_out_s <= color_out_d;
		end if;
	end process;
	 
end Behavioral;