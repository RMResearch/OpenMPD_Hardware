library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity PinMapping is
	port (
		clk		   : in  std_logic;
		address_in  : in  std_logic_vector (7 downto 0);
		address_out : out std_logic_vector (7 downto 0)
	);
end PinMapping;

architecture Behavioral of PinMapping is
	
	signal address_out_s	: std_logic_vector (7 downto 0) := (others => '0');
	signal address_out_d	: std_logic_vector (7 downto 0) := (others => '0');

	subtype PIN is std_logic_vector(7 downto 0);
	type ROM is array (0 to 255) of PIN;
	constant pin_ROM : ROM := (
	"11111001", "11111101", "11110001", "11110101", "11101001", "11101101", "11100001", "11100101", "11011001", "11011101", "11010001", "11010101", "11001001", "11001101", "11000001", "11000101",
	"11111000", "11111100", "11110000", "11110100", "11101000", "11101100", "11100000", "11100100", "11011000", "11011100", "11010000", "11010100", "11001000", "11001100", "11000000", "11000100",
	"11111011", "11111110", "11110011", "11110110", "11101011", "11101110", "11100011", "11100110", "11011011", "11011110", "11010011", "11010110", "11001011", "11001110", "11000011", "11000110",
	"11111010", "11111111", "11110010", "11110111", "11101010", "11101111", "11100010", "11100111", "11011010", "11011111", "11010010", "11010111", "11001010", "11001111", "11000010", "11000111",
	"10111001", "10111101", "10110001", "10110101", "10101001", "10101101", "10100001", "10100101", "10011001", "10011101", "10010001", "10010101", "10001001", "10001101", "10000001", "10000101",
	"10111000", "10111100", "10110000", "10110100", "10101000", "10101100", "10100000", "10100100", "10011000", "10011100", "10010000", "10010100", "10001000", "10001100", "10000000", "10000100",
	"10111011", "10111110", "10110011", "10110110", "10101011", "10101110", "10100011", "10100110", "10011011", "10011110", "10010011", "10010110", "10001011", "10001110", "10000011", "10000110",
	"10111010", "10111111", "10110010", "10110111", "10101010", "10101111", "10100010", "10100111", "10011010", "10011111", "10010010", "10010111", "10001010", "10001111", "10000010", "10000111",
	"01111001", "01111101", "01110001", "01110101", "01101001", "01101101", "01100001", "01100101", "01011001", "01011101", "01010001", "01010101", "01001001", "01001101", "01000001", "01000101",
	"01111000", "01111100", "01110000", "01110100", "01101000", "01101100", "01100000", "01100100", "01011000", "01011100", "01010000", "01010100", "01001000", "01001100", "01000000", "01000100",
	"01111011", "01111110", "01110011", "01110110", "01101011", "01101110", "01100011", "01100110", "01011011", "01011110", "01010011", "01010110", "01001011", "01001110", "01000011", "01000110",
	"01111010", "01111111", "01110010", "01110111", "01101010", "01101111", "01100010", "01100111", "01011010", "01011111", "01010010", "01010111", "01001010", "01001111", "01000010", "01000111",
	"00111001", "00111101", "00110001", "00110101", "00101001", "00101101", "00100001", "00100101", "00011001", "00011101", "00010001", "00010101", "00001001", "00001101", "00000001", "00000101",
	"00111000", "00111100", "00110000", "00110100", "00101000", "00101100", "00100000", "00100100", "00011000", "00011100", "00010000", "00010100", "00001000", "00001100", "00000000", "00000100",
	"00111011", "00111110", "00110011", "00110110", "00101011", "00101110", "00100011", "00100110", "00011011", "00011110", "00010011", "00010110", "00001011", "00001110", "00000011", "00000110",
	"00111010", "00111111", "00110010", "00110111", "00101010", "00101111", "00100010", "00100111", "00011010", "00011111", "00010010", "00010111", "00001010", "00001111", "00000010", "00000111"

--		"11000101","11000100","11000110","11000111","10000101","10000100","10000110","10000111","01000101","01000100","01000110","01000111","00000101","00000100","00000110","00000111",
--		"11000001","11000000","11000011","11000010","10000001","10000000","10000011","10000010","01000001","01000000","01000011","01000010","00000001","00000000","00000011","00000010",
--		"11001101","11001100","11001110","11001111","10001101","10001100","10001110","10001111","01001101","01001100","01001110","01001111","00001101","00001100","00001110","00001111",
--		"11001001","11001000","11001011","11001010","10001001","10001000","10001011","10001010","01001001","01001000","01001011","01001010","00001001","00001000","00001011","00001010",
--		"11010101","11010100","11010110","11010111","10010101","10010100","10010110","10010111","01010101","01010100","01010110","01010111","00010101","00010100","00010110","00010111",
--		"11010001","11010000","11010011","11010010","10010001","10010000","10010011","10010010","01010001","01010000","01010011","01010010","00010001","00010000","00010011","00010010",
--		"11011101","11011100","11011110","11011111","10011101","10011100","10011110","10011111","01011101","01011100","01011110","01011111","00011101","00011100","00011110","00011111",
--		"11011001","11011000","11011011","11011010","10011001","10011000","10011011","10011010","01011001","01011000","01011011","01011010","00011001","00011000","00011011","00011010",
--		"11100101","11100100","11100110","11100111","10100101","10100100","10100110","10100111","01100101","01100100","01100110","01100111","00100101","00100100","00100110","00100111",
--		"11100001","11100000","11100011","11100010","10100001","10100000","10100011","10100010","01100001","01100000","01100011","01100010","00100001","00100000","00100011","00100010",
--		"11101101","11101100","11101110","11101111","10101101","10101100","10101110","10101111","01101101","01101100","01101110","01101111","00101101","00101100","00101110","00101111",
--		"11101001","11101000","11101011","11101010","10101001","10101000","10101011","10101010","01101001","01101000","01101011","01101010","00101001","00101000","00101011","00101010",
--		"11110101","11110100","11110110","11110111","10110101","10110100","10110110","10110111","01110101","01110100","01110110","01110111","00110101","00110100","00110110","00110111",
--		"11110001","11110000","11110011","11110010","10110001","10110000","10110011","10110010","01110001","01110000","01110011","01110010","00110001","00110000","00110011","00110010",
--		"11111101","11111100","11111110","11111111","10111101","10111100","10111110","10111111","01111101","01111100","01111110","01111111","00111101","00111100","00111110","00111111",
--		"11111001","11111000","11111011","11111010","10111001","10111000","10111011","10111010","01111001","01111000","01111011","01111010","00111001","00111000","00111011","00111010"
	);	
	
begin
	
	address_out <= address_out_s;
	
	process (clk) begin
		if rising_edge(clk) then
			address_out_d <= address_in;--pin_ROM(CONV_INTEGER(address_in));
			address_out_s <= address_out_d;
		end if;
	end process;
end Behavioral;