AmplitudeCorrectionLUT_inst : AmplitudeCorrectionLUT PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
